module mux_for (
	input 			i0 , 
	input 			i1 , 
	input 			i2 , 
	input 			i3 , 
	input 	[1:0] 		sel, 
	output 	 	reg	y
);


wire [3:0] i_int;
assign i_int = {i3,i2,i1,i0};
integer k;

always @ (*)
	begin
	y = 0;
	for(k = 0; k < 4; k=k+1) begin
		if(k == sel)
			y = i_int[k];
	end
end

endmodule


