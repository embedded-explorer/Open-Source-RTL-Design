module sub_module(
	input 	a , 
	input 	b , 
	output 	y
);
 	assign y = a & b;
endmodule


module multiple_module_opt2(
	input 	a , 
	input 	b , 
	input 	c , 
	input 	d , 
	output 	y
);

wire n1,n2,n3;

sub_module U1 (.a(a)	, .b(1'b0)	, .y(n1));
sub_module U2 (.a(b)	, .b(c) 	, .y(n2));
sub_module U3 (.a(n2)	, .b(d) 	, .y(n3));
sub_module U4 (.a(n3)	, .b(n1) 	, .y(y)	);

endmodule
