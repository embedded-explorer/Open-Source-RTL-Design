module sub_module1(
	input 	a , 
	input 	b , 
	output	y
);
 	assign y = a & b;
endmodule


module sub_module2(
	input 	a , 
	input 	b , 
	output 	y
);
 	assign y = a^b;
endmodule


module multiple_module_opt1(
	input 	a , 
	input 	b , 
	input 	c , 
	input 	d , 
	output 	y	
);

wire n1,n2,n3;

sub_module1 U1 (.a(a)	, .b(1'b1) 	, .y(n1));
sub_module2 U2 (.a(n1)	, .b(1'b0) 	, .y(n2));
sub_module2 U3 (.a(b)	, .b(d) 	, .y(n3));

assign y = c | (b & n1); 

endmodule
