module rca (
	input 	[7:0] 	num1 , 
	input 	[7:0] 	num2 , 
	output 	[8:0] 	sum
);	

wire 	[7:0] 	int_sum;
wire 	[7:0]	int_co;

genvar i;
generate
	for (i = 1 ; i < 8; i=i+1) begin
		fa u_fa_1 (.a(num1[i]),.b(num2[i]),.c(int_co[i-1]),.co(int_co[i]),.sum(int_sum[i]));
	end

endgenerate

fa u_fa_0 (
	.a(num1[0]),
	.b(num2[0]),
	.c(1'b0),
	.co(int_co[0]),
	.sum(int_sum[0])
	);


assign sum[7:0] = int_sum;
assign sum[8] = int_co[7];

endmodule

