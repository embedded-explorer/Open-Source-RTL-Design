module counter_opt1 (
	input 	clk , 
	input 	reset , 
	output 	q
);

reg [2:0] count;

assign q = count[0];

always @(posedge clk ,posedge reset)
begin
	if(reset)
		count <= 3'b000;
	else
		count <= count + 1;
end

endmodule
