module counter_opt2 (
	input 	clk , 
	input 	reset , 
	output 	q
);

reg [2:0] count;

assign q = (count[2:0] == 3'b100);

always @(posedge clk ,posedge reset)
begin
	if(reset)
		count <= 3'b000;
	else
		count <= count + 1;
end

endmodule
