module bad_mux (
	input 		i0 , 
	input 		i1 , 
	input 		sel, 
	output 	reg 	y
);

always @ (sel)
begin
	if(sel)
		y <= i1;
	else 
		y <= i0;
end

endmodule
