module fa (
	input 	a , 
	input 	b , 
	input 	c , 
	output 	co, 
	output 	sum
);
	assign {co,sum}  = a + b + c ;
endmodule
