module demux_case (
	output 		o0 , 
	output 		o1 , 
	output 		o2 , 
	output 		o3 , 
	output 		o4 , 
	output 		o5 , 
	output 		o6 , 
	output 		o7 , 
	input 	[2:0] 	sel  , 
	input 		i
);

reg [7:0]y_int;
assign {o7,o6,o5,o4,o3,o2,o1,o0} = y_int;
integer k;

always @ (*)
begin
y_int = 8'b0;
	case(sel)
		3'b000 : y_int[0] = i;
		3'b001 : y_int[1] = i;
		3'b010 : y_int[2] = i;
		3'b011 : y_int[3] = i;
		3'b100 : y_int[4] = i;
		3'b101 : y_int[5] = i;
		3'b110 : y_int[6] = i;
		3'b111 : y_int[7] = i;
	endcase

end

endmodule


