module dff_const1(
	input 		clk, 
	input 		reset, 
	output 	reg 	q
);

always @(posedge clk, posedge reset)
begin
	if(reset)
		q <= 1'b0;
	else
		q <= 1'b1;
end

endmodule
